`ifndef _CMPTYPES_H_
`define _CMPTYPES_H_

localparam EQ = 3'b000;
localparam NE = 3'b001;
localparam LT = 3'b010;
localparam LE = 3'b011;
localparam GE = 3'b100;
localparam GT = 3'b101;

`endif